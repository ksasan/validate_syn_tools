module m;

initial
  $display("Hello World");
endmodule
